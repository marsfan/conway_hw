--- Testbench for POPCOUNT_ARITH

-- This Source Code Form is subject to the terms of the Mozilla Public
-- License, v. 2.0. If a copy of the MPL was not distributed with this
-- file, You can obtain one at https://mozilla.org/MPL/2.0/.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library vunit_lib;
context vunit_lib.vunit_context;

entity POPCOUNT_ARITH_TB is
    generic (
        runner_cfg : string
    );
end entity POPCOUNT_ARITH_TB;

architecture TEST of POPCOUNT_ARITH_TB is

    component POPCOUNT_ARITH is
        port (
            N     : in  std_logic;
            NE    : in  std_logic;
            E     : in  std_logic;
            SE    : in  std_logic;
            S     : in  std_logic;
            SW    : in  std_logic;
            W     : in  std_logic;
            NW    : in  std_logic;
            COUNT : out std_logic_vector(3 downto 0)
        );
    end component POPCOUNT_ARITH;

    -- Array of test cases to evaluate

    type test_record is record
        N     : std_logic;
        NE    : std_logic;
        E     : std_logic;
        SE    : std_logic;
        S     : std_logic;
        SW    : std_logic;
        W     : std_logic;
        NW    : std_logic;
        COUNT : std_logic_vector(3 downto 0);
    end record test_record;

    type test_array_t is array (natural range <>) of test_record;

    constant TEST_ARRAY : test_array_t := (
        ('0', '0', '0', '0', '0', '0', '0', '0', "0000"),
        ('0', '0', '0', '0', '0', '0', '0', '1', "0001"),
        ('0', '0', '0', '0', '0', '0', '1', '0', "0001"),
        ('0', '0', '0', '0', '0', '0', '1', '1', "0010"),
        ('0', '0', '0', '0', '0', '1', '0', '0', "0001"),
        ('0', '0', '0', '0', '0', '1', '0', '1', "0010"),
        ('0', '0', '0', '0', '0', '1', '1', '0', "0010"),
        ('0', '0', '0', '0', '0', '1', '1', '1', "0011"),
        ('0', '0', '0', '0', '1', '0', '0', '0', "0001"),
        ('0', '0', '0', '0', '1', '0', '0', '1', "0010"),
        ('0', '0', '0', '0', '1', '0', '1', '0', "0010"),
        ('0', '0', '0', '0', '1', '0', '1', '1', "0011"),
        ('0', '0', '0', '0', '1', '1', '0', '0', "0010"),
        ('0', '0', '0', '0', '1', '1', '0', '1', "0011"),
        ('0', '0', '0', '0', '1', '1', '1', '0', "0011"),
        ('0', '0', '0', '0', '1', '1', '1', '1', "0100"),
        ('0', '0', '0', '1', '0', '0', '0', '0', "0001"),
        ('0', '0', '0', '1', '0', '0', '0', '1', "0010"),
        ('0', '0', '0', '1', '0', '0', '1', '0', "0010"),
        ('0', '0', '0', '1', '0', '0', '1', '1', "0011"),
        ('0', '0', '0', '1', '0', '1', '0', '0', "0010"),
        ('0', '0', '0', '1', '0', '1', '0', '1', "0011"),
        ('0', '0', '0', '1', '0', '1', '1', '0', "0011"),
        ('0', '0', '0', '1', '0', '1', '1', '1', "0100"),
        ('0', '0', '0', '1', '1', '0', '0', '0', "0010"),
        ('0', '0', '0', '1', '1', '0', '0', '1', "0011"),
        ('0', '0', '0', '1', '1', '0', '1', '0', "0011"),
        ('0', '0', '0', '1', '1', '0', '1', '1', "0100"),
        ('0', '0', '0', '1', '1', '1', '0', '0', "0011"),
        ('0', '0', '0', '1', '1', '1', '0', '1', "0100"),
        ('0', '0', '0', '1', '1', '1', '1', '0', "0100"),
        ('0', '0', '0', '1', '1', '1', '1', '1', "0101"),
        ('0', '0', '1', '0', '0', '0', '0', '0', "0001"),
        ('0', '0', '1', '0', '0', '0', '0', '1', "0010"),
        ('0', '0', '1', '0', '0', '0', '1', '0', "0010"),
        ('0', '0', '1', '0', '0', '0', '1', '1', "0011"),
        ('0', '0', '1', '0', '0', '1', '0', '0', "0010"),
        ('0', '0', '1', '0', '0', '1', '0', '1', "0011"),
        ('0', '0', '1', '0', '0', '1', '1', '0', "0011"),
        ('0', '0', '1', '0', '0', '1', '1', '1', "0100"),
        ('0', '0', '1', '0', '1', '0', '0', '0', "0010"),
        ('0', '0', '1', '0', '1', '0', '0', '1', "0011"),
        ('0', '0', '1', '0', '1', '0', '1', '0', "0011"),
        ('0', '0', '1', '0', '1', '0', '1', '1', "0100"),
        ('0', '0', '1', '0', '1', '1', '0', '0', "0011"),
        ('0', '0', '1', '0', '1', '1', '0', '1', "0100"),
        ('0', '0', '1', '0', '1', '1', '1', '0', "0100"),
        ('0', '0', '1', '0', '1', '1', '1', '1', "0101"),
        ('0', '0', '1', '1', '0', '0', '0', '0', "0010"),
        ('0', '0', '1', '1', '0', '0', '0', '1', "0011"),
        ('0', '0', '1', '1', '0', '0', '1', '0', "0011"),
        ('0', '0', '1', '1', '0', '0', '1', '1', "0100"),
        ('0', '0', '1', '1', '0', '1', '0', '0', "0011"),
        ('0', '0', '1', '1', '0', '1', '0', '1', "0100"),
        ('0', '0', '1', '1', '0', '1', '1', '0', "0100"),
        ('0', '0', '1', '1', '0', '1', '1', '1', "0101"),
        ('0', '0', '1', '1', '1', '0', '0', '0', "0011"),
        ('0', '0', '1', '1', '1', '0', '0', '1', "0100"),
        ('0', '0', '1', '1', '1', '0', '1', '0', "0100"),
        ('0', '0', '1', '1', '1', '0', '1', '1', "0101"),
        ('0', '0', '1', '1', '1', '1', '0', '0', "0100"),
        ('0', '0', '1', '1', '1', '1', '0', '1', "0101"),
        ('0', '0', '1', '1', '1', '1', '1', '0', "0101"),
        ('0', '0', '1', '1', '1', '1', '1', '1', "0110"),
        ('0', '1', '0', '0', '0', '0', '0', '0', "0001"),
        ('0', '1', '0', '0', '0', '0', '0', '1', "0010"),
        ('0', '1', '0', '0', '0', '0', '1', '0', "0010"),
        ('0', '1', '0', '0', '0', '0', '1', '1', "0011"),
        ('0', '1', '0', '0', '0', '1', '0', '0', "0010"),
        ('0', '1', '0', '0', '0', '1', '0', '1', "0011"),
        ('0', '1', '0', '0', '0', '1', '1', '0', "0011"),
        ('0', '1', '0', '0', '0', '1', '1', '1', "0100"),
        ('0', '1', '0', '0', '1', '0', '0', '0', "0010"),
        ('0', '1', '0', '0', '1', '0', '0', '1', "0011"),
        ('0', '1', '0', '0', '1', '0', '1', '0', "0011"),
        ('0', '1', '0', '0', '1', '0', '1', '1', "0100"),
        ('0', '1', '0', '0', '1', '1', '0', '0', "0011"),
        ('0', '1', '0', '0', '1', '1', '0', '1', "0100"),
        ('0', '1', '0', '0', '1', '1', '1', '0', "0100"),
        ('0', '1', '0', '0', '1', '1', '1', '1', "0101"),
        ('0', '1', '0', '1', '0', '0', '0', '0', "0010"),
        ('0', '1', '0', '1', '0', '0', '0', '1', "0011"),
        ('0', '1', '0', '1', '0', '0', '1', '0', "0011"),
        ('0', '1', '0', '1', '0', '0', '1', '1', "0100"),
        ('0', '1', '0', '1', '0', '1', '0', '0', "0011"),
        ('0', '1', '0', '1', '0', '1', '0', '1', "0100"),
        ('0', '1', '0', '1', '0', '1', '1', '0', "0100"),
        ('0', '1', '0', '1', '0', '1', '1', '1', "0101"),
        ('0', '1', '0', '1', '1', '0', '0', '0', "0011"),
        ('0', '1', '0', '1', '1', '0', '0', '1', "0100"),
        ('0', '1', '0', '1', '1', '0', '1', '0', "0100"),
        ('0', '1', '0', '1', '1', '0', '1', '1', "0101"),
        ('0', '1', '0', '1', '1', '1', '0', '0', "0100"),
        ('0', '1', '0', '1', '1', '1', '0', '1', "0101"),
        ('0', '1', '0', '1', '1', '1', '1', '0', "0101"),
        ('0', '1', '0', '1', '1', '1', '1', '1', "0110"),
        ('0', '1', '1', '0', '0', '0', '0', '0', "0010"),
        ('0', '1', '1', '0', '0', '0', '0', '1', "0011"),
        ('0', '1', '1', '0', '0', '0', '1', '0', "0011"),
        ('0', '1', '1', '0', '0', '0', '1', '1', "0100"),
        ('0', '1', '1', '0', '0', '1', '0', '0', "0011"),
        ('0', '1', '1', '0', '0', '1', '0', '1', "0100"),
        ('0', '1', '1', '0', '0', '1', '1', '0', "0100"),
        ('0', '1', '1', '0', '0', '1', '1', '1', "0101"),
        ('0', '1', '1', '0', '1', '0', '0', '0', "0011"),
        ('0', '1', '1', '0', '1', '0', '0', '1', "0100"),
        ('0', '1', '1', '0', '1', '0', '1', '0', "0100"),
        ('0', '1', '1', '0', '1', '0', '1', '1', "0101"),
        ('0', '1', '1', '0', '1', '1', '0', '0', "0100"),
        ('0', '1', '1', '0', '1', '1', '0', '1', "0101"),
        ('0', '1', '1', '0', '1', '1', '1', '0', "0101"),
        ('0', '1', '1', '0', '1', '1', '1', '1', "0110"),
        ('0', '1', '1', '1', '0', '0', '0', '0', "0011"),
        ('0', '1', '1', '1', '0', '0', '0', '1', "0100"),
        ('0', '1', '1', '1', '0', '0', '1', '0', "0100"),
        ('0', '1', '1', '1', '0', '0', '1', '1', "0101"),
        ('0', '1', '1', '1', '0', '1', '0', '0', "0100"),
        ('0', '1', '1', '1', '0', '1', '0', '1', "0101"),
        ('0', '1', '1', '1', '0', '1', '1', '0', "0101"),
        ('0', '1', '1', '1', '0', '1', '1', '1', "0110"),
        ('0', '1', '1', '1', '1', '0', '0', '0', "0100"),
        ('0', '1', '1', '1', '1', '0', '0', '1', "0101"),
        ('0', '1', '1', '1', '1', '0', '1', '0', "0101"),
        ('0', '1', '1', '1', '1', '0', '1', '1', "0110"),
        ('0', '1', '1', '1', '1', '1', '0', '0', "0101"),
        ('0', '1', '1', '1', '1', '1', '0', '1', "0110"),
        ('0', '1', '1', '1', '1', '1', '1', '0', "0110"),
        ('0', '1', '1', '1', '1', '1', '1', '1', "0111"),
        ('1', '0', '0', '0', '0', '0', '0', '0', "0001"),
        ('1', '0', '0', '0', '0', '0', '0', '1', "0010"),
        ('1', '0', '0', '0', '0', '0', '1', '0', "0010"),
        ('1', '0', '0', '0', '0', '0', '1', '1', "0011"),
        ('1', '0', '0', '0', '0', '1', '0', '0', "0010"),
        ('1', '0', '0', '0', '0', '1', '0', '1', "0011"),
        ('1', '0', '0', '0', '0', '1', '1', '0', "0011"),
        ('1', '0', '0', '0', '0', '1', '1', '1', "0100"),
        ('1', '0', '0', '0', '1', '0', '0', '0', "0010"),
        ('1', '0', '0', '0', '1', '0', '0', '1', "0011"),
        ('1', '0', '0', '0', '1', '0', '1', '0', "0011"),
        ('1', '0', '0', '0', '1', '0', '1', '1', "0100"),
        ('1', '0', '0', '0', '1', '1', '0', '0', "0011"),
        ('1', '0', '0', '0', '1', '1', '0', '1', "0100"),
        ('1', '0', '0', '0', '1', '1', '1', '0', "0100"),
        ('1', '0', '0', '0', '1', '1', '1', '1', "0101"),
        ('1', '0', '0', '1', '0', '0', '0', '0', "0010"),
        ('1', '0', '0', '1', '0', '0', '0', '1', "0011"),
        ('1', '0', '0', '1', '0', '0', '1', '0', "0011"),
        ('1', '0', '0', '1', '0', '0', '1', '1', "0100"),
        ('1', '0', '0', '1', '0', '1', '0', '0', "0011"),
        ('1', '0', '0', '1', '0', '1', '0', '1', "0100"),
        ('1', '0', '0', '1', '0', '1', '1', '0', "0100"),
        ('1', '0', '0', '1', '0', '1', '1', '1', "0101"),
        ('1', '0', '0', '1', '1', '0', '0', '0', "0011"),
        ('1', '0', '0', '1', '1', '0', '0', '1', "0100"),
        ('1', '0', '0', '1', '1', '0', '1', '0', "0100"),
        ('1', '0', '0', '1', '1', '0', '1', '1', "0101"),
        ('1', '0', '0', '1', '1', '1', '0', '0', "0100"),
        ('1', '0', '0', '1', '1', '1', '0', '1', "0101"),
        ('1', '0', '0', '1', '1', '1', '1', '0', "0101"),
        ('1', '0', '0', '1', '1', '1', '1', '1', "0110"),
        ('1', '0', '1', '0', '0', '0', '0', '0', "0010"),
        ('1', '0', '1', '0', '0', '0', '0', '1', "0011"),
        ('1', '0', '1', '0', '0', '0', '1', '0', "0011"),
        ('1', '0', '1', '0', '0', '0', '1', '1', "0100"),
        ('1', '0', '1', '0', '0', '1', '0', '0', "0011"),
        ('1', '0', '1', '0', '0', '1', '0', '1', "0100"),
        ('1', '0', '1', '0', '0', '1', '1', '0', "0100"),
        ('1', '0', '1', '0', '0', '1', '1', '1', "0101"),
        ('1', '0', '1', '0', '1', '0', '0', '0', "0011"),
        ('1', '0', '1', '0', '1', '0', '0', '1', "0100"),
        ('1', '0', '1', '0', '1', '0', '1', '0', "0100"),
        ('1', '0', '1', '0', '1', '0', '1', '1', "0101"),
        ('1', '0', '1', '0', '1', '1', '0', '0', "0100"),
        ('1', '0', '1', '0', '1', '1', '0', '1', "0101"),
        ('1', '0', '1', '0', '1', '1', '1', '0', "0101"),
        ('1', '0', '1', '0', '1', '1', '1', '1', "0110"),
        ('1', '0', '1', '1', '0', '0', '0', '0', "0011"),
        ('1', '0', '1', '1', '0', '0', '0', '1', "0100"),
        ('1', '0', '1', '1', '0', '0', '1', '0', "0100"),
        ('1', '0', '1', '1', '0', '0', '1', '1', "0101"),
        ('1', '0', '1', '1', '0', '1', '0', '0', "0100"),
        ('1', '0', '1', '1', '0', '1', '0', '1', "0101"),
        ('1', '0', '1', '1', '0', '1', '1', '0', "0101"),
        ('1', '0', '1', '1', '0', '1', '1', '1', "0110"),
        ('1', '0', '1', '1', '1', '0', '0', '0', "0100"),
        ('1', '0', '1', '1', '1', '0', '0', '1', "0101"),
        ('1', '0', '1', '1', '1', '0', '1', '0', "0101"),
        ('1', '0', '1', '1', '1', '0', '1', '1', "0110"),
        ('1', '0', '1', '1', '1', '1', '0', '0', "0101"),
        ('1', '0', '1', '1', '1', '1', '0', '1', "0110"),
        ('1', '0', '1', '1', '1', '1', '1', '0', "0110"),
        ('1', '0', '1', '1', '1', '1', '1', '1', "0111"),
        ('1', '1', '0', '0', '0', '0', '0', '0', "0010"),
        ('1', '1', '0', '0', '0', '0', '0', '1', "0011"),
        ('1', '1', '0', '0', '0', '0', '1', '0', "0011"),
        ('1', '1', '0', '0', '0', '0', '1', '1', "0100"),
        ('1', '1', '0', '0', '0', '1', '0', '0', "0011"),
        ('1', '1', '0', '0', '0', '1', '0', '1', "0100"),
        ('1', '1', '0', '0', '0', '1', '1', '0', "0100"),
        ('1', '1', '0', '0', '0', '1', '1', '1', "0101"),
        ('1', '1', '0', '0', '1', '0', '0', '0', "0011"),
        ('1', '1', '0', '0', '1', '0', '0', '1', "0100"),
        ('1', '1', '0', '0', '1', '0', '1', '0', "0100"),
        ('1', '1', '0', '0', '1', '0', '1', '1', "0101"),
        ('1', '1', '0', '0', '1', '1', '0', '0', "0100"),
        ('1', '1', '0', '0', '1', '1', '0', '1', "0101"),
        ('1', '1', '0', '0', '1', '1', '1', '0', "0101"),
        ('1', '1', '0', '0', '1', '1', '1', '1', "0110"),
        ('1', '1', '0', '1', '0', '0', '0', '0', "0011"),
        ('1', '1', '0', '1', '0', '0', '0', '1', "0100"),
        ('1', '1', '0', '1', '0', '0', '1', '0', "0100"),
        ('1', '1', '0', '1', '0', '0', '1', '1', "0101"),
        ('1', '1', '0', '1', '0', '1', '0', '0', "0100"),
        ('1', '1', '0', '1', '0', '1', '0', '1', "0101"),
        ('1', '1', '0', '1', '0', '1', '1', '0', "0101"),
        ('1', '1', '0', '1', '0', '1', '1', '1', "0110"),
        ('1', '1', '0', '1', '1', '0', '0', '0', "0100"),
        ('1', '1', '0', '1', '1', '0', '0', '1', "0101"),
        ('1', '1', '0', '1', '1', '0', '1', '0', "0101"),
        ('1', '1', '0', '1', '1', '0', '1', '1', "0110"),
        ('1', '1', '0', '1', '1', '1', '0', '0', "0101"),
        ('1', '1', '0', '1', '1', '1', '0', '1', "0110"),
        ('1', '1', '0', '1', '1', '1', '1', '0', "0110"),
        ('1', '1', '0', '1', '1', '1', '1', '1', "0111"),
        ('1', '1', '1', '0', '0', '0', '0', '0', "0011"),
        ('1', '1', '1', '0', '0', '0', '0', '1', "0100"),
        ('1', '1', '1', '0', '0', '0', '1', '0', "0100"),
        ('1', '1', '1', '0', '0', '0', '1', '1', "0101"),
        ('1', '1', '1', '0', '0', '1', '0', '0', "0100"),
        ('1', '1', '1', '0', '0', '1', '0', '1', "0101"),
        ('1', '1', '1', '0', '0', '1', '1', '0', "0101"),
        ('1', '1', '1', '0', '0', '1', '1', '1', "0110"),
        ('1', '1', '1', '0', '1', '0', '0', '0', "0100"),
        ('1', '1', '1', '0', '1', '0', '0', '1', "0101"),
        ('1', '1', '1', '0', '1', '0', '1', '0', "0101"),
        ('1', '1', '1', '0', '1', '0', '1', '1', "0110"),
        ('1', '1', '1', '0', '1', '1', '0', '0', "0101"),
        ('1', '1', '1', '0', '1', '1', '0', '1', "0110"),
        ('1', '1', '1', '0', '1', '1', '1', '0', "0110"),
        ('1', '1', '1', '0', '1', '1', '1', '1', "0111"),
        ('1', '1', '1', '1', '0', '0', '0', '0', "0100"),
        ('1', '1', '1', '1', '0', '0', '0', '1', "0101"),
        ('1', '1', '1', '1', '0', '0', '1', '0', "0101"),
        ('1', '1', '1', '1', '0', '0', '1', '1', "0110"),
        ('1', '1', '1', '1', '0', '1', '0', '0', "0101"),
        ('1', '1', '1', '1', '0', '1', '0', '1', "0110"),
        ('1', '1', '1', '1', '0', '1', '1', '0', "0110"),
        ('1', '1', '1', '1', '0', '1', '1', '1', "0111"),
        ('1', '1', '1', '1', '1', '0', '0', '0', "0101"),
        ('1', '1', '1', '1', '1', '0', '0', '1', "0110"),
        ('1', '1', '1', '1', '1', '0', '1', '0', "0110"),
        ('1', '1', '1', '1', '1', '0', '1', '1', "0111"),
        ('1', '1', '1', '1', '1', '1', '0', '0', "0110"),
        ('1', '1', '1', '1', '1', '1', '0', '1', "0111"),
        ('1', '1', '1', '1', '1', '1', '1', '0', "0111"),
        ('1', '1', '1', '1', '1', '1', '1', '1', "1000")
    );

    signal N     : std_logic;
    signal NE    : std_logic;
    signal E     : std_logic;
    signal SE    : std_logic;
    signal S     : std_logic;
    signal SW    : std_logic;
    signal W     : std_logic;
    signal NW    : std_logic;
    signal COUNT : std_logic_vector(3 downto 0);

begin

    test_popcount : POPCOUNT_ARITH
        port map (
            N     => N,
            NE    => NE,
            E     => E,
            SE    => SE,
            S     => S,
            SW    => SW,
            W     => W,
            NW    => NW,
            COUNT => COUNT
        );

    test_proc : process is
    begin

        test_runner_setup(runner, runner_cfg);

        if run("TEST_POPCOUNT_ARITH") then

            for i in TEST_ARRAY'range loop

                -- Set all signal
                N  <= TEST_ARRAY(i).N;
                NE <= TEST_ARRAY(i).NE;
                E  <= TEST_ARRAY(i).E;
                SE <= TEST_ARRAY(i).SE;
                S  <= TEST_ARRAY(i).S;
                SW <= TEST_ARRAY(i).SW;
                W  <= TEST_ARRAY(i).W;
                NW <= TEST_ARRAY(i).NW;

                wait for 1 ns;
                -- Check output
                check_equal(COUNT, TEST_ARRAY(i).COUNT, "COUNT");

            end loop;

        end if;

        test_runner_cleanup(runner);

    end process test_proc;

end architecture TEST;
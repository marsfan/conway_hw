/*
 * Copyright (c) 2024 Your Name
 * SPDX-License-Identifier: Apache-2.0
 */

`default_nettype none

/* svlint off keyword_forbidden_wire_reg */
module tt_um_conway (
    input  wire [7:0] ui_in,    // Dedicated inputs
    output wire [7:0] uo_out,   // Dedicated outputs
    input  wire [7:0] uio_in,   // IOs: Input path
    output wire [7:0] uio_out,  // IOs: Output path
    output wire [7:0] uio_oe,   // IOs: Enable path (active high: 0=input, 1=output)
    input  wire       ena,      // always 1 when the design is powered, so you can ignore it
    input  wire       clk,      // clock
    input  wire       rst_n     // reset_n - low to reset
);
  /* svlint on keyword_forbidden_wire_reg */

  conway_8x8_serial_v4 conway_mod(
    .data_in(ui_in[0]),
    .mode(ui_in[2:1]),
    .reset(rst_n),
    .clk(clk),
    .data_out(uo_out[0]),
    .din_led(uo_out[1]),
    .clk_led(uo_out[2]),
    .dout_led(uo_out[3]),
    .mode_leds(uo_out[5:4])
  );

  // All output pins must be assigned. If not used, assign to 0.
  // assign uo_out  = ui_in + uio_in;  // Example: ou_out is the sum of ui_in and uio_in
  assign uio_out = 0;
  assign uio_oe  = 0;

  assign uo_out[7:6] = 0;

  // List all unused inputs to prevent warnings

endmodule

--- Testbench for POPCOUNT_ARITH

-- This Source Code Form is subject to the terms of the Mozilla Public
-- License, v. 2.0. If a copy of the MPL was not distributed with this
-- file, You can obtain one at https: //mozilla.org/MPL/2.0/.
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library vunit_lib;
context vunit_lib.vunit_context;

entity POPCOUNT_ARITH_TB is
    generic (runner_cfg : string);
end entity POPCOUNT_ARITH_TB;

architecture TEST of POPCOUNT_ARITH_TB is

    component POPCOUNT_ARITH is
        port (
            N     : in std_logic;
            NE    : in std_logic;
            E     : in std_logic;
            SE    : in std_logic;
            S     : in std_logic;
            SW    : in std_logic;
            W     : in std_logic;
            NW    : in std_logic;
            COUNT : out std_logic_vector(3 downto 0)
        );
    end component POPCOUNT_ARITH;

    --- Array of test cases to evaluate
    type test_record is record
        -- Inputs
        N     : std_logic;
        NE    : std_logic;
        E     : std_logic;
        SE    : std_logic;
        S     : std_logic;
        SW    : std_logic;
        W     : std_logic;
        NW    : std_logic;

        -- outputs
        COUNT : std_logic_vector(3 downto 0);
    end record;
    type test_array_t is array (natural range <>) of test_record;
    constant test_array : test_array_t := (
        ('0', '0', '0', '0', '0', '0', '0', '0', "0000"),
        ('0', '0', '0', '0', '0', '0', '0', '1', "0001"),
        ('0', '0', '0', '0', '0', '0', '1', '0', "0001"),
        ('0', '0', '0', '0', '0', '0', '1', '1', "0010"),
        ('0', '0', '0', '0', '0', '1', '0', '0', "0001"),
        ('0', '0', '0', '0', '0', '1', '0', '1', "0010"),
        ('0', '0', '0', '0', '0', '1', '1', '0', "0010"),
        ('0', '0', '0', '0', '0', '1', '1', '1', "0011"),
        ('0', '0', '0', '0', '1', '0', '0', '0', "0001"),
        ('0', '0', '0', '0', '1', '0', '0', '1', "0010"),
        ('0', '0', '0', '0', '1', '0', '1', '0', "0010"),
        ('0', '0', '0', '0', '1', '0', '1', '1', "0011"),
        ('0', '0', '0', '0', '1', '1', '0', '0', "0010"),
        ('0', '0', '0', '0', '1', '1', '0', '1', "0011"),
        ('0', '0', '0', '0', '1', '1', '1', '0', "0011"),
        ('0', '0', '0', '0', '1', '1', '1', '1', "0100"),
        ('0', '0', '0', '1', '0', '0', '0', '0', "0001"),
        ('0', '0', '0', '1', '0', '0', '0', '1', "0010"),
        ('0', '0', '0', '1', '0', '0', '1', '0', "0010"),
        ('0', '0', '0', '1', '0', '0', '1', '1', "0011"),
        ('0', '0', '0', '1', '0', '1', '0', '0', "0010"),
        ('0', '0', '0', '1', '0', '1', '0', '1', "0011"),
        ('0', '0', '0', '1', '0', '1', '1', '0', "0011"),
        ('0', '0', '0', '1', '0', '1', '1', '1', "0100"),
        ('0', '0', '0', '1', '1', '0', '0', '0', "0010"),
        ('0', '0', '0', '1', '1', '0', '0', '1', "0011"),
        ('0', '0', '0', '1', '1', '0', '1', '0', "0011"),
        ('0', '0', '0', '1', '1', '0', '1', '1', "0100"),
        ('0', '0', '0', '1', '1', '1', '0', '0', "0011"),
        ('0', '0', '0', '1', '1', '1', '0', '1', "0100"),
        ('0', '0', '0', '1', '1', '1', '1', '0', "0100"),
        ('0', '0', '0', '1', '1', '1', '1', '1', "0101"),
        ('0', '0', '1', '0', '0', '0', '0', '0', "0001"),
        ('0', '0', '1', '0', '0', '0', '0', '1', "0010"),
        ('0', '0', '1', '0', '0', '0', '1', '0', "0010"),
        ('0', '0', '1', '0', '0', '0', '1', '1', "0011"),
        ('0', '0', '1', '0', '0', '1', '0', '0', "0010"),
        ('0', '0', '1', '0', '0', '1', '0', '1', "0011"),
        ('0', '0', '1', '0', '0', '1', '1', '0', "0011"),
        ('0', '0', '1', '0', '0', '1', '1', '1', "0100"),
        ('0', '0', '1', '0', '1', '0', '0', '0', "0010"),
        ('0', '0', '1', '0', '1', '0', '0', '1', "0011"),
        ('0', '0', '1', '0', '1', '0', '1', '0', "0011"),
        ('0', '0', '1', '0', '1', '0', '1', '1', "0100"),
        ('0', '0', '1', '0', '1', '1', '0', '0', "0011"),
        ('0', '0', '1', '0', '1', '1', '0', '1', "0100"),
        ('0', '0', '1', '0', '1', '1', '1', '0', "0100"),
        ('0', '0', '1', '0', '1', '1', '1', '1', "0101"),
        ('0', '0', '1', '1', '0', '0', '0', '0', "0010"),
        ('0', '0', '1', '1', '0', '0', '0', '1', "0011"),
        ('0', '0', '1', '1', '0', '0', '1', '0', "0011"),
        ('0', '0', '1', '1', '0', '0', '1', '1', "0100"),
        ('0', '0', '1', '1', '0', '1', '0', '0', "0011"),
        ('0', '0', '1', '1', '0', '1', '0', '1', "0100"),
        ('0', '0', '1', '1', '0', '1', '1', '0', "0100"),
        ('0', '0', '1', '1', '0', '1', '1', '1', "0101"),
        ('0', '0', '1', '1', '1', '0', '0', '0', "0011"),
        ('0', '0', '1', '1', '1', '0', '0', '1', "0100"),
        ('0', '0', '1', '1', '1', '0', '1', '0', "0100"),
        ('0', '0', '1', '1', '1', '0', '1', '1', "0101"),
        ('0', '0', '1', '1', '1', '1', '0', '0', "0100"),
        ('0', '0', '1', '1', '1', '1', '0', '1', "0101"),
        ('0', '0', '1', '1', '1', '1', '1', '0', "0101"),
        ('0', '0', '1', '1', '1', '1', '1', '1', "0110"),
        ('0', '1', '0', '0', '0', '0', '0', '0', "0001"),
        ('0', '1', '0', '0', '0', '0', '0', '1', "0010"),
        ('0', '1', '0', '0', '0', '0', '1', '0', "0010"),
        ('0', '1', '0', '0', '0', '0', '1', '1', "0011"),
        ('0', '1', '0', '0', '0', '1', '0', '0', "0010"),
        ('0', '1', '0', '0', '0', '1', '0', '1', "0011"),
        ('0', '1', '0', '0', '0', '1', '1', '0', "0011"),
        ('0', '1', '0', '0', '0', '1', '1', '1', "0100"),
        ('0', '1', '0', '0', '1', '0', '0', '0', "0010"),
        ('0', '1', '0', '0', '1', '0', '0', '1', "0011"),
        ('0', '1', '0', '0', '1', '0', '1', '0', "0011"),
        ('0', '1', '0', '0', '1', '0', '1', '1', "0100"),
        ('0', '1', '0', '0', '1', '1', '0', '0', "0011"),
        ('0', '1', '0', '0', '1', '1', '0', '1', "0100"),
        ('0', '1', '0', '0', '1', '1', '1', '0', "0100"),
        ('0', '1', '0', '0', '1', '1', '1', '1', "0101"),
        ('0', '1', '0', '1', '0', '0', '0', '0', "0010"),
        ('0', '1', '0', '1', '0', '0', '0', '1', "0011"),
        ('0', '1', '0', '1', '0', '0', '1', '0', "0011"),
        ('0', '1', '0', '1', '0', '0', '1', '1', "0100"),
        ('0', '1', '0', '1', '0', '1', '0', '0', "0011"),
        ('0', '1', '0', '1', '0', '1', '0', '1', "0100"),
        ('0', '1', '0', '1', '0', '1', '1', '0', "0100"),
        ('0', '1', '0', '1', '0', '1', '1', '1', "0101"),
        ('0', '1', '0', '1', '1', '0', '0', '0', "0011"),
        ('0', '1', '0', '1', '1', '0', '0', '1', "0100"),
        ('0', '1', '0', '1', '1', '0', '1', '0', "0100"),
        ('0', '1', '0', '1', '1', '0', '1', '1', "0101"),
        ('0', '1', '0', '1', '1', '1', '0', '0', "0100"),
        ('0', '1', '0', '1', '1', '1', '0', '1', "0101"),
        ('0', '1', '0', '1', '1', '1', '1', '0', "0101"),
        ('0', '1', '0', '1', '1', '1', '1', '1', "0110"),
        ('0', '1', '1', '0', '0', '0', '0', '0', "0010"),
        ('0', '1', '1', '0', '0', '0', '0', '1', "0011"),
        ('0', '1', '1', '0', '0', '0', '1', '0', "0011"),
        ('0', '1', '1', '0', '0', '0', '1', '1', "0100"),
        ('0', '1', '1', '0', '0', '1', '0', '0', "0011"),
        ('0', '1', '1', '0', '0', '1', '0', '1', "0100"),
        ('0', '1', '1', '0', '0', '1', '1', '0', "0100"),
        ('0', '1', '1', '0', '0', '1', '1', '1', "0101"),
        ('0', '1', '1', '0', '1', '0', '0', '0', "0011"),
        ('0', '1', '1', '0', '1', '0', '0', '1', "0100"),
        ('0', '1', '1', '0', '1', '0', '1', '0', "0100"),
        ('0', '1', '1', '0', '1', '0', '1', '1', "0101"),
        ('0', '1', '1', '0', '1', '1', '0', '0', "0100"),
        ('0', '1', '1', '0', '1', '1', '0', '1', "0101"),
        ('0', '1', '1', '0', '1', '1', '1', '0', "0101"),
        ('0', '1', '1', '0', '1', '1', '1', '1', "0110"),
        ('0', '1', '1', '1', '0', '0', '0', '0', "0011"),
        ('0', '1', '1', '1', '0', '0', '0', '1', "0100"),
        ('0', '1', '1', '1', '0', '0', '1', '0', "0100"),
        ('0', '1', '1', '1', '0', '0', '1', '1', "0101"),
        ('0', '1', '1', '1', '0', '1', '0', '0', "0100"),
        ('0', '1', '1', '1', '0', '1', '0', '1', "0101"),
        ('0', '1', '1', '1', '0', '1', '1', '0', "0101"),
        ('0', '1', '1', '1', '0', '1', '1', '1', "0110"),
        ('0', '1', '1', '1', '1', '0', '0', '0', "0100"),
        ('0', '1', '1', '1', '1', '0', '0', '1', "0101"),
        ('0', '1', '1', '1', '1', '0', '1', '0', "0101"),
        ('0', '1', '1', '1', '1', '0', '1', '1', "0110"),
        ('0', '1', '1', '1', '1', '1', '0', '0', "0101"),
        ('0', '1', '1', '1', '1', '1', '0', '1', "0110"),
        ('0', '1', '1', '1', '1', '1', '1', '0', "0110"),
        ('0', '1', '1', '1', '1', '1', '1', '1', "0111"),
        ('1', '0', '0', '0', '0', '0', '0', '0', "0001"),
        ('1', '0', '0', '0', '0', '0', '0', '1', "0010"),
        ('1', '0', '0', '0', '0', '0', '1', '0', "0010"),
        ('1', '0', '0', '0', '0', '0', '1', '1', "0011"),
        ('1', '0', '0', '0', '0', '1', '0', '0', "0010"),
        ('1', '0', '0', '0', '0', '1', '0', '1', "0011"),
        ('1', '0', '0', '0', '0', '1', '1', '0', "0011"),
        ('1', '0', '0', '0', '0', '1', '1', '1', "0100"),
        ('1', '0', '0', '0', '1', '0', '0', '0', "0010"),
        ('1', '0', '0', '0', '1', '0', '0', '1', "0011"),
        ('1', '0', '0', '0', '1', '0', '1', '0', "0011"),
        ('1', '0', '0', '0', '1', '0', '1', '1', "0100"),
        ('1', '0', '0', '0', '1', '1', '0', '0', "0011"),
        ('1', '0', '0', '0', '1', '1', '0', '1', "0100"),
        ('1', '0', '0', '0', '1', '1', '1', '0', "0100"),
        ('1', '0', '0', '0', '1', '1', '1', '1', "0101"),
        ('1', '0', '0', '1', '0', '0', '0', '0', "0010"),
        ('1', '0', '0', '1', '0', '0', '0', '1', "0011"),
        ('1', '0', '0', '1', '0', '0', '1', '0', "0011"),
        ('1', '0', '0', '1', '0', '0', '1', '1', "0100"),
        ('1', '0', '0', '1', '0', '1', '0', '0', "0011"),
        ('1', '0', '0', '1', '0', '1', '0', '1', "0100"),
        ('1', '0', '0', '1', '0', '1', '1', '0', "0100"),
        ('1', '0', '0', '1', '0', '1', '1', '1', "0101"),
        ('1', '0', '0', '1', '1', '0', '0', '0', "0011"),
        ('1', '0', '0', '1', '1', '0', '0', '1', "0100"),
        ('1', '0', '0', '1', '1', '0', '1', '0', "0100"),
        ('1', '0', '0', '1', '1', '0', '1', '1', "0101"),
        ('1', '0', '0', '1', '1', '1', '0', '0', "0100"),
        ('1', '0', '0', '1', '1', '1', '0', '1', "0101"),
        ('1', '0', '0', '1', '1', '1', '1', '0', "0101"),
        ('1', '0', '0', '1', '1', '1', '1', '1', "0110"),
        ('1', '0', '1', '0', '0', '0', '0', '0', "0010"),
        ('1', '0', '1', '0', '0', '0', '0', '1', "0011"),
        ('1', '0', '1', '0', '0', '0', '1', '0', "0011"),
        ('1', '0', '1', '0', '0', '0', '1', '1', "0100"),
        ('1', '0', '1', '0', '0', '1', '0', '0', "0011"),
        ('1', '0', '1', '0', '0', '1', '0', '1', "0100"),
        ('1', '0', '1', '0', '0', '1', '1', '0', "0100"),
        ('1', '0', '1', '0', '0', '1', '1', '1', "0101"),
        ('1', '0', '1', '0', '1', '0', '0', '0', "0011"),
        ('1', '0', '1', '0', '1', '0', '0', '1', "0100"),
        ('1', '0', '1', '0', '1', '0', '1', '0', "0100"),
        ('1', '0', '1', '0', '1', '0', '1', '1', "0101"),
        ('1', '0', '1', '0', '1', '1', '0', '0', "0100"),
        ('1', '0', '1', '0', '1', '1', '0', '1', "0101"),
        ('1', '0', '1', '0', '1', '1', '1', '0', "0101"),
        ('1', '0', '1', '0', '1', '1', '1', '1', "0110"),
        ('1', '0', '1', '1', '0', '0', '0', '0', "0011"),
        ('1', '0', '1', '1', '0', '0', '0', '1', "0100"),
        ('1', '0', '1', '1', '0', '0', '1', '0', "0100"),
        ('1', '0', '1', '1', '0', '0', '1', '1', "0101"),
        ('1', '0', '1', '1', '0', '1', '0', '0', "0100"),
        ('1', '0', '1', '1', '0', '1', '0', '1', "0101"),
        ('1', '0', '1', '1', '0', '1', '1', '0', "0101"),
        ('1', '0', '1', '1', '0', '1', '1', '1', "0110"),
        ('1', '0', '1', '1', '1', '0', '0', '0', "0100"),
        ('1', '0', '1', '1', '1', '0', '0', '1', "0101"),
        ('1', '0', '1', '1', '1', '0', '1', '0', "0101"),
        ('1', '0', '1', '1', '1', '0', '1', '1', "0110"),
        ('1', '0', '1', '1', '1', '1', '0', '0', "0101"),
        ('1', '0', '1', '1', '1', '1', '0', '1', "0110"),
        ('1', '0', '1', '1', '1', '1', '1', '0', "0110"),
        ('1', '0', '1', '1', '1', '1', '1', '1', "0111"),
        ('1', '1', '0', '0', '0', '0', '0', '0', "0010"),
        ('1', '1', '0', '0', '0', '0', '0', '1', "0011"),
        ('1', '1', '0', '0', '0', '0', '1', '0', "0011"),
        ('1', '1', '0', '0', '0', '0', '1', '1', "0100"),
        ('1', '1', '0', '0', '0', '1', '0', '0', "0011"),
        ('1', '1', '0', '0', '0', '1', '0', '1', "0100"),
        ('1', '1', '0', '0', '0', '1', '1', '0', "0100"),
        ('1', '1', '0', '0', '0', '1', '1', '1', "0101"),
        ('1', '1', '0', '0', '1', '0', '0', '0', "0011"),
        ('1', '1', '0', '0', '1', '0', '0', '1', "0100"),
        ('1', '1', '0', '0', '1', '0', '1', '0', "0100"),
        ('1', '1', '0', '0', '1', '0', '1', '1', "0101"),
        ('1', '1', '0', '0', '1', '1', '0', '0', "0100"),
        ('1', '1', '0', '0', '1', '1', '0', '1', "0101"),
        ('1', '1', '0', '0', '1', '1', '1', '0', "0101"),
        ('1', '1', '0', '0', '1', '1', '1', '1', "0110"),
        ('1', '1', '0', '1', '0', '0', '0', '0', "0011"),
        ('1', '1', '0', '1', '0', '0', '0', '1', "0100"),
        ('1', '1', '0', '1', '0', '0', '1', '0', "0100"),
        ('1', '1', '0', '1', '0', '0', '1', '1', "0101"),
        ('1', '1', '0', '1', '0', '1', '0', '0', "0100"),
        ('1', '1', '0', '1', '0', '1', '0', '1', "0101"),
        ('1', '1', '0', '1', '0', '1', '1', '0', "0101"),
        ('1', '1', '0', '1', '0', '1', '1', '1', "0110"),
        ('1', '1', '0', '1', '1', '0', '0', '0', "0100"),
        ('1', '1', '0', '1', '1', '0', '0', '1', "0101"),
        ('1', '1', '0', '1', '1', '0', '1', '0', "0101"),
        ('1', '1', '0', '1', '1', '0', '1', '1', "0110"),
        ('1', '1', '0', '1', '1', '1', '0', '0', "0101"),
        ('1', '1', '0', '1', '1', '1', '0', '1', "0110"),
        ('1', '1', '0', '1', '1', '1', '1', '0', "0110"),
        ('1', '1', '0', '1', '1', '1', '1', '1', "0111"),
        ('1', '1', '1', '0', '0', '0', '0', '0', "0011"),
        ('1', '1', '1', '0', '0', '0', '0', '1', "0100"),
        ('1', '1', '1', '0', '0', '0', '1', '0', "0100"),
        ('1', '1', '1', '0', '0', '0', '1', '1', "0101"),
        ('1', '1', '1', '0', '0', '1', '0', '0', "0100"),
        ('1', '1', '1', '0', '0', '1', '0', '1', "0101"),
        ('1', '1', '1', '0', '0', '1', '1', '0', "0101"),
        ('1', '1', '1', '0', '0', '1', '1', '1', "0110"),
        ('1', '1', '1', '0', '1', '0', '0', '0', "0100"),
        ('1', '1', '1', '0', '1', '0', '0', '1', "0101"),
        ('1', '1', '1', '0', '1', '0', '1', '0', "0101"),
        ('1', '1', '1', '0', '1', '0', '1', '1', "0110"),
        ('1', '1', '1', '0', '1', '1', '0', '0', "0101"),
        ('1', '1', '1', '0', '1', '1', '0', '1', "0110"),
        ('1', '1', '1', '0', '1', '1', '1', '0', "0110"),
        ('1', '1', '1', '0', '1', '1', '1', '1', "0111"),
        ('1', '1', '1', '1', '0', '0', '0', '0', "0100"),
        ('1', '1', '1', '1', '0', '0', '0', '1', "0101"),
        ('1', '1', '1', '1', '0', '0', '1', '0', "0101"),
        ('1', '1', '1', '1', '0', '0', '1', '1', "0110"),
        ('1', '1', '1', '1', '0', '1', '0', '0', "0101"),
        ('1', '1', '1', '1', '0', '1', '0', '1', "0110"),
        ('1', '1', '1', '1', '0', '1', '1', '0', "0110"),
        ('1', '1', '1', '1', '0', '1', '1', '1', "0111"),
        ('1', '1', '1', '1', '1', '0', '0', '0', "0101"),
        ('1', '1', '1', '1', '1', '0', '0', '1', "0110"),
        ('1', '1', '1', '1', '1', '0', '1', '0', "0110"),
        ('1', '1', '1', '1', '1', '0', '1', '1', "0111"),
        ('1', '1', '1', '1', '1', '1', '0', '0', "0110"),
        ('1', '1', '1', '1', '1', '1', '0', '1', "0111"),
        ('1', '1', '1', '1', '1', '1', '1', '0', "0111"),
        ('1', '1', '1', '1', '1', '1', '1', '1', "1000")
    );

    signal  N, NE, E, SE, S, SW, W, NW : std_logic;
    signal COUNT : std_logic_vector(3 downto 0);

begin

    TEST_POPCOUNT : POPCOUNT_ARITH port map(
        N =>  N,
        NE =>  NE,
        E =>  E,
        SE =>  SE,
        S =>  S,
        SW =>  SW,
        W =>  W,
        NW =>  NW,
        COUNT =>  COUNT
    );

    test_proc : process
    begin
        test_runner_setup(runner, runner_cfg);
        if run("TEST_POPCOUNT_ARITH") then
            for i in test_array'range loop
                -- Set all signal
                N <= test_array(i).N;
                NE <= test_array(i).NE;
                E <= test_array(i).E;
                SE <= test_array(i).SE;
                S <= test_array(i).S;
                SW <= test_array(i).SW;
                W <= test_array(i).W;
                NW <= test_array(i).NW;

                wait for 1 ns;
                -- Check output
                check_equal(COUNT, test_array(i).COUNT, "COUNT");
            end loop;
        end if;
        test_runner_cleanup(runner);

    end process;

end architecture;
/*
* This Source Code Form is subject to the terms of the Mozilla Public
* License, v. 2.0. If a copy of the MPL was not distributed with this
* file, You can obtain one at https: //mozilla.org/MPL/2.0/.
*/

`include "tests/test_utils.sv"

module cell_grid_tb();

    logic [63:0] INPUT_STATE;
    logic [63:0] NEXT_STATE;

    CELL_GRID #(8, 8) dut (
        .INPUT_STATE(INPUT_STATE),
        .NEXT_STATE(NEXT_STATE)
    );

    initial begin
        int errcount;
        errcount = 0;

        // Configure to dump variables to VCD file
        $dumpfile("waveforms/cell_grid_tb.vcd");
        $dumpvars(0, cell_grid_tb);

        // Testing a few of the different patterns from the
        // Wikipedia page on conway's game of life.

        INPUT_STATE <= 64'h0000001818000000;
        #1
        `CHECK_EQ(NEXT_STATE, 64'h0000001818000000, errcount, "Block");

        INPUT_STATE <= 64'h0000102828100000;
        #1
        `CHECK_EQ(NEXT_STATE, 64'h0000102828100000, errcount, "Behive");

        INPUT_STATE <= 64'h0000001010100000;
        #1
        `CHECK_EQ(NEXT_STATE, 64'h0000000038000000, errcount, "Blinker");

        INPUT_STATE <= 64'h0060601818000000;
        #1
        `CHECK_EQ(NEXT_STATE, 64'h0060400818000000, errcount, "Beacon");

        INPUT_STATE <= 64'hC080000000000000;
        #1
        `CHECK_EQ(NEXT_STATE, 64'hC0C0000000000000, errcount, "Corner1");

        INPUT_STATE <= 64'h8080800000000000;
        #1
        `CHECK_EQ(NEXT_STATE, 64'h00C0000000000000, errcount, "Corner2");

        `STOP_IF_ERR(errcount);


    end

endmodule